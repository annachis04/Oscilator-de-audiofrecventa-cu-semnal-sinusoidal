LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY SCHEMATIC1 IS 

END SCHEMATIC1;



ARCHITECTURE STRUCTURE OF SCHEMATIC1 IS

-- COMPONENTS

COMPONENT \1k\
	PORT (
	\2\ : INOUT std_logic;
	\1\ : INOUT std_logic
	); END COMPONENT;

COMPONENT \50k\
	PORT (
	\2\ : INOUT std_logic;
	\1\ : INOUT std_logic;
	t : INOUT std_logic
	); END COMPONENT;

COMPONENT QBC846B
	PORT (
	B : IN std_logic;
	E : INOUT std_logic;
	C : INOUT std_logic
	); END COMPONENT;

COMPONENT QBC856B
	PORT (
	B : IN std_logic;
	E : INOUT std_logic;
	C : INOUT std_logic
	); END COMPONENT;

COMPONENT QBC846B
	PORT (
	B : IN std_logic;
	E : INOUT std_logic;
	C : INOUT std_logic
	); END COMPONENT;

COMPONENT QBC846B
	PORT (
	B : IN std_logic;
	E : INOUT std_logic;
	C : INOUT std_logic
	); END COMPONENT;

COMPONENT \V-\
	PORT (
	\1\ : INOUT std_logic
	); END COMPONENT;

COMPONENT \33n\
	PORT (
	\1\ : INOUT std_logic;
	\2\ : INOUT std_logic
	); END COMPONENT;

COMPONENT CON2
	PORT (
	\1\ : INOUT std_logic;
	\2\ : INOUT std_logic
	); END COMPONENT;

COMPONENT D1N4148
	PORT (
	\1\ : INOUT std_logic;
	\2\ : INOUT std_logic
	); END COMPONENT;

COMPONENT D1N4148
	PORT (
	\1\ : INOUT std_logic;
	\2\ : INOUT std_logic
	); END COMPONENT;

COMPONENT \5V,LED,LED\
	PORT (
	\1\ : INOUT std_logic;
	\2\ : INOUT std_logic
	); END COMPONENT;

COMPONENT QBC856B
	PORT (
	B : IN std_logic;
	E : INOUT std_logic;
	C : INOUT std_logic
	); END COMPONENT;

COMPONENT QBC856B
	PORT (
	B : IN std_logic;
	E : INOUT std_logic;
	C : INOUT std_logic
	); END COMPONENT;

COMPONENT QBC846B
	PORT (
	B : IN std_logic;
	E : INOUT std_logic;
	C : INOUT std_logic
	); END COMPONENT;

-- SIGNALS

SIGNAL GND : std_logic;
SIGNAL N97649 : std_logic;
SIGNAL N977031 : std_logic;
SIGNAL N977231 : std_logic;
SIGNAL N97755 : std_logic;
SIGNAL N97835 : std_logic;
SIGNAL N97875 : std_logic;
SIGNAL N97939 : std_logic;
SIGNAL N97965 : std_logic;
SIGNAL N97969 : std_logic;
SIGNAL N97983 : std_logic;
SIGNAL N98131 : std_logic;
SIGNAL N98141 : std_logic;
SIGNAL N98201 : std_logic;
SIGNAL N98233 : std_logic;
SIGNAL N983391 : std_logic;
SIGNAL N98425 : std_logic;
SIGNAL N98451 : std_logic;
SIGNAL N98621 : std_logic;
SIGNAL N98633 : std_logic;
SIGNAL N98691 : std_logic;

-- INSTANCE ATTRIBUTES

ATTRIBUTE SLOPE:string;
ATTRIBUTE SLOPE of R25 : label is "RSMAX";
ATTRIBUTE TC2:string;
ATTRIBUTE TC2 of R25 : label is "0";
ATTRIBUTE TC1:string;
ATTRIBUTE TC1 of R25 : label is "0";
ATTRIBUTE MAX_TEMP:string;
ATTRIBUTE MAX_TEMP of R25 : label is "RTMAX";
ATTRIBUTE DIST:string;
ATTRIBUTE DIST of R25 : label is "FLAT";
ATTRIBUTE VOLTAGE:string;
ATTRIBUTE VOLTAGE of R25 : label is "RVMAX";
ATTRIBUTE POWER:string;
ATTRIBUTE POWER of R25 : label is "RMAX";
ATTRIBUTE PSPICETEMPLATE:string;
ATTRIBUTE PSPICETEMPLATE of R25 : label is "R^@REFDES %1 %2 ?TOLERANCE|R^@REFDES| @VALUE TC=@TC1,@TC2 ?TOLERANCE|\n.model R^@REFDES RES R=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2|";
ATTRIBUTE SLOPE of R26 : label is "RSMAX";
ATTRIBUTE TC2 of R26 : label is "0";
ATTRIBUTE TC1 of R26 : label is "0";
ATTRIBUTE MAX_TEMP of R26 : label is "RTMAX";
ATTRIBUTE DIST of R26 : label is "FLAT";
ATTRIBUTE VOLTAGE of R26 : label is "RVMAX";
ATTRIBUTE POWER of R26 : label is "RMAX";
ATTRIBUTE PSPICETEMPLATE of R26 : label is "R^@REFDES %1 %2 ?TOLERANCE|R^@REFDES| @VALUE TC=@TC1,@TC2 ?TOLERANCE|\n.model R^@REFDES RES R=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2|";
ATTRIBUTE SET:string;
ATTRIBUTE SET of R27 : label is "0.1";
ATTRIBUTE PSPICETEMPLATE of R27 : label is "X^@REFDES %1 %T %2 POT PARAMS: SET=@SET VALUE=@VALUE";
ATTRIBUTE SET of R28 : label is "0.1";
ATTRIBUTE PSPICETEMPLATE of R28 : label is "X^@REFDES %1 %T %2 POT PARAMS: SET=@SET VALUE=@VALUE";
ATTRIBUTE SLOPE of R29 : label is "RSMAX";
ATTRIBUTE TC2 of R29 : label is "0";
ATTRIBUTE TC1 of R29 : label is "0";
ATTRIBUTE MAX_TEMP of R29 : label is "RTMAX";
ATTRIBUTE DIST of R29 : label is "FLAT";
ATTRIBUTE VOLTAGE of R29 : label is "RVMAX";
ATTRIBUTE POWER of R29 : label is "RMAX";
ATTRIBUTE PSPICETEMPLATE of R29 : label is "R^@REFDES %1 %2 ?TOLERANCE|R^@REFDES| @VALUE TC=@TC1,@TC2 ?TOLERANCE|\n.model R^@REFDES RES R=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2|";
ATTRIBUTE PSPICETEMPLATE of Q20 : label is "Q^@REFDES %C %B %E @MODEL ?AREA/@AREA/";
ATTRIBUTE PSPICETEMPLATE of Q21 : label is "Q^@REFDES %C %B %E @MODEL ?AREA/@AREA/";
ATTRIBUTE PSPICETEMPLATE of Q22 : label is "Q^@REFDES %C %B %E @MODEL ?AREA/@AREA/";
ATTRIBUTE PSPICETEMPLATE of Q23 : label is "Q^@REFDES %C %B %E @MODEL ?AREA/@AREA/";
ATTRIBUTE SLOPE of R30 : label is "RSMAX";
ATTRIBUTE TC2 of R30 : label is "0";
ATTRIBUTE TC1 of R30 : label is "0";
ATTRIBUTE MAX_TEMP of R30 : label is "RTMAX";
ATTRIBUTE DIST of R30 : label is "FLAT";
ATTRIBUTE VOLTAGE of R30 : label is "RVMAX";
ATTRIBUTE POWER of R30 : label is "RMAX";
ATTRIBUTE PSPICETEMPLATE of R30 : label is "R^@REFDES %1 %2 ?TOLERANCE|R^@REFDES| @VALUE TC=@TC1,@TC2 ?TOLERANCE|\n.model R^@REFDES RES R=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2|";
ATTRIBUTE SLOPE of R31 : label is "RSMAX";
ATTRIBUTE TC2 of R31 : label is "0";
ATTRIBUTE TC1 of R31 : label is "0";
ATTRIBUTE MAX_TEMP of R31 : label is "RTMAX";
ATTRIBUTE DIST of R31 : label is "FLAT";
ATTRIBUTE VOLTAGE of R31 : label is "RVMAX";
ATTRIBUTE POWER of R31 : label is "RMAX";
ATTRIBUTE PSPICETEMPLATE of R31 : label is "R^@REFDES %1 %2 ?TOLERANCE|R^@REFDES| @VALUE TC=@TC1,@TC2 ?TOLERANCE|\n.model R^@REFDES RES R=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2|";
ATTRIBUTE SET of R32 : label is "0.1";
ATTRIBUTE PSPICETEMPLATE of R32 : label is "X^@REFDES %1 %T %2 POT PARAMS: SET=@SET VALUE=@VALUE";
ATTRIBUTE SLOPE of R33 : label is "RSMAX";
ATTRIBUTE TC2 of R33 : label is "0";
ATTRIBUTE TC1 of R33 : label is "0";
ATTRIBUTE MAX_TEMP of R33 : label is "RTMAX";
ATTRIBUTE DIST of R33 : label is "FLAT";
ATTRIBUTE VOLTAGE of R33 : label is "RVMAX";
ATTRIBUTE POWER of R33 : label is "RMAX";
ATTRIBUTE PSPICETEMPLATE of R33 : label is "R^@REFDES %1 %2 ?TOLERANCE|R^@REFDES| @VALUE TC=@TC1,@TC2 ?TOLERANCE|\n.model R^@REFDES RES R=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2|";
ATTRIBUTE SLOPE of R7 : label is "RSMAX";
ATTRIBUTE TC2 of R7 : label is "0";
ATTRIBUTE TC1 of R7 : label is "0";
ATTRIBUTE MAX_TEMP of R7 : label is "RTMAX";
ATTRIBUTE DIST of R7 : label is "FLAT";
ATTRIBUTE VOLTAGE of R7 : label is "RVMAX";
ATTRIBUTE POWER of R7 : label is "RMAX";
ATTRIBUTE PSPICETEMPLATE of R7 : label is "R^@REFDES %1 %2 ?TOLERANCE|R^@REFDES| @VALUE TC=@TC1,@TC2 ?TOLERANCE|\n.model R^@REFDES RES R=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2|";
ATTRIBUTE SLOPE of R8 : label is "RSMAX";
ATTRIBUTE TC2 of R8 : label is "0";
ATTRIBUTE TC1 of R8 : label is "0";
ATTRIBUTE MAX_TEMP of R8 : label is "RTMAX";
ATTRIBUTE DIST of R8 : label is "FLAT";
ATTRIBUTE VOLTAGE of R8 : label is "RVMAX";
ATTRIBUTE POWER of R8 : label is "RMAX";
ATTRIBUTE PSPICETEMPLATE of R8 : label is "R^@REFDES %1 %2 ?TOLERANCE|R^@REFDES| @VALUE TC=@TC1,@TC2 ?TOLERANCE|\n.model R^@REFDES RES R=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2|";
ATTRIBUTE SLOPE of C6 : label is "CSMAX";
ATTRIBUTE KNEE:string;
ATTRIBUTE KNEE of C6 : label is "CBMAX";
ATTRIBUTE TC2 of C6 : label is "0";
ATTRIBUTE CURRENT:string;
ATTRIBUTE CURRENT of C6 : label is "CIMAX";
ATTRIBUTE VC1:string;
ATTRIBUTE VC1 of C6 : label is "0";
ATTRIBUTE VC2:string;
ATTRIBUTE VC2 of C6 : label is "0";
ATTRIBUTE MAX_TEMP of C6 : label is "CTMAX";
ATTRIBUTE DIST of C6 : label is "FLAT";
ATTRIBUTE TC1 of C6 : label is "0";
ATTRIBUTE VOLTAGE of C6 : label is "CMAX";
ATTRIBUTE PSPICETEMPLATE of C6 : label is "C^@REFDES %1 %2 ?TOLERANCE|C^@REFDES| @VALUE ?IC/IC=@IC/ TC=@TC1,@TC2 ?TOLERANCE|\n.model C^@REFDES CAP C=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2 VC1=@VC1 VC2=@VC2|";
ATTRIBUTE SLOPE of C7 : label is "CSMAX";
ATTRIBUTE KNEE of C7 : label is "CBMAX";
ATTRIBUTE TC2 of C7 : label is "0";
ATTRIBUTE CURRENT of C7 : label is "CIMAX";
ATTRIBUTE VC1 of C7 : label is "0";
ATTRIBUTE VC2 of C7 : label is "0";
ATTRIBUTE MAX_TEMP of C7 : label is "CTMAX";
ATTRIBUTE DIST of C7 : label is "FLAT";
ATTRIBUTE TC1 of C7 : label is "0";
ATTRIBUTE VOLTAGE of C7 : label is "CMAX";
ATTRIBUTE PSPICETEMPLATE of C7 : label is "C^@REFDES %1 %2 ?TOLERANCE|C^@REFDES| @VALUE ?IC/IC=@IC/ TC=@TC1,@TC2 ?TOLERANCE|\n.model C^@REFDES CAP C=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2 VC1=@VC1 VC2=@VC2|";
ATTRIBUTE SLOPE of C8 : label is "CSMAX";
ATTRIBUTE KNEE of C8 : label is "CBMAX";
ATTRIBUTE TC2 of C8 : label is "0";
ATTRIBUTE CURRENT of C8 : label is "CIMAX";
ATTRIBUTE VC1 of C8 : label is "0";
ATTRIBUTE VC2 of C8 : label is "0";
ATTRIBUTE MAX_TEMP of C8 : label is "CTMAX";
ATTRIBUTE DIST of C8 : label is "FLAT";
ATTRIBUTE TC1 of C8 : label is "0";
ATTRIBUTE VOLTAGE of C8 : label is "CMAX";
ATTRIBUTE PSPICETEMPLATE of C8 : label is "C^@REFDES %1 %2 ?TOLERANCE|C^@REFDES| @VALUE ?IC/IC=@IC/ TC=@TC1,@TC2 ?TOLERANCE|\n.model C^@REFDES CAP C=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2 VC1=@VC1 VC2=@VC2|";
ATTRIBUTE \COMPONENT\:string;
ATTRIBUTE \COMPONENT\ of D1 : label is "1N4148";
ATTRIBUTE PSPICETEMPLATE of D1 : label is "D^@REFDES %1 %2 @MODEL ?AREA/@AREA/";
ATTRIBUTE SLOPE of R19 : label is "RSMAX";
ATTRIBUTE TC2 of R19 : label is "0";
ATTRIBUTE TC1 of R19 : label is "0";
ATTRIBUTE MAX_TEMP of R19 : label is "RTMAX";
ATTRIBUTE DIST of R19 : label is "FLAT";
ATTRIBUTE VOLTAGE of R19 : label is "RVMAX";
ATTRIBUTE POWER of R19 : label is "RMAX";
ATTRIBUTE PSPICETEMPLATE of R19 : label is "R^@REFDES %1 %2 ?TOLERANCE|R^@REFDES| @VALUE TC=@TC1,@TC2 ?TOLERANCE|\n.model R^@REFDES RES R=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2|";
ATTRIBUTE \COMPONENT\ of D2 : label is "1N4148";
ATTRIBUTE PSPICETEMPLATE of D2 : label is "D^@REFDES %1 %2 @MODEL ?AREA/@AREA/";
ATTRIBUTE \IS\:string;
ATTRIBUTE \IS\ of D3 : label is "1.7603e-027";
ATTRIBUTE VR:string;
ATTRIBUTE VR of D3 : label is "5";
ATTRIBUTE PSPICEMODELINGAPPTYPE:string;
ATTRIBUTE PSPICEMODELINGAPPTYPE of D3 : label is "LED";
ATTRIBUTE BV:string;
ATTRIBUTE BV of D3 : label is "5";
ATTRIBUTE \IF\:string;
ATTRIBUTE \IF\ of D3 : label is "30E-3";
ATTRIBUTE PDM:string;
ATTRIBUTE PDM of D3 : label is "114E-3";
ATTRIBUTE IBV:string;
ATTRIBUTE IBV of D3 : label is "5e-6";
ATTRIBUTE APPPROP:string;
ATTRIBUTE APPPROP of D3 : label is "mN=LED,fV=3,fC=20E-3";
ATTRIBUTE RS:string;
ATTRIBUTE RS of D3 : label is "2";
ATTRIBUTE PSPICETEMPLATE of Q17 : label is "Q^@REFDES %C %B %E @MODEL ?AREA/@AREA/";
ATTRIBUTE PSPICETEMPLATE of Q18 : label is "Q^@REFDES %C %B %E @MODEL ?AREA/@AREA/";
ATTRIBUTE PSPICETEMPLATE of Q19 : label is "Q^@REFDES %C %B %E @MODEL ?AREA/@AREA/";
ATTRIBUTE SLOPE of R20 : label is "RSMAX";
ATTRIBUTE TC2 of R20 : label is "0";
ATTRIBUTE TC1 of R20 : label is "0";
ATTRIBUTE MAX_TEMP of R20 : label is "RTMAX";
ATTRIBUTE DIST of R20 : label is "FLAT";
ATTRIBUTE VOLTAGE of R20 : label is "RVMAX";
ATTRIBUTE POWER of R20 : label is "RMAX";
ATTRIBUTE PSPICETEMPLATE of R20 : label is "R^@REFDES %1 %2 ?TOLERANCE|R^@REFDES| @VALUE TC=@TC1,@TC2 ?TOLERANCE|\n.model R^@REFDES RES R=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2|";
ATTRIBUTE SLOPE of R22 : label is "RSMAX";
ATTRIBUTE TC2 of R22 : label is "0";
ATTRIBUTE TC1 of R22 : label is "0";
ATTRIBUTE MAX_TEMP of R22 : label is "RTMAX";
ATTRIBUTE DIST of R22 : label is "FLAT";
ATTRIBUTE VOLTAGE of R22 : label is "RVMAX";
ATTRIBUTE POWER of R22 : label is "RMAX";
ATTRIBUTE PSPICETEMPLATE of R22 : label is "R^@REFDES %1 %2 ?TOLERANCE|R^@REFDES| @VALUE TC=@TC1,@TC2 ?TOLERANCE|\n.model R^@REFDES RES R=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2|";
ATTRIBUTE SLOPE of R23 : label is "RSMAX";
ATTRIBUTE TC2 of R23 : label is "0";
ATTRIBUTE TC1 of R23 : label is "0";
ATTRIBUTE MAX_TEMP of R23 : label is "RTMAX";
ATTRIBUTE DIST of R23 : label is "FLAT";
ATTRIBUTE VOLTAGE of R23 : label is "RVMAX";
ATTRIBUTE POWER of R23 : label is "RMAX";
ATTRIBUTE PSPICETEMPLATE of R23 : label is "R^@REFDES %1 %2 ?TOLERANCE|R^@REFDES| @VALUE TC=@TC1,@TC2 ?TOLERANCE|\n.model R^@REFDES RES R=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2|";
ATTRIBUTE SLOPE of R24 : label is "RSMAX";
ATTRIBUTE TC2 of R24 : label is "0";
ATTRIBUTE TC1 of R24 : label is "0";
ATTRIBUTE MAX_TEMP of R24 : label is "RTMAX";
ATTRIBUTE DIST of R24 : label is "FLAT";
ATTRIBUTE VOLTAGE of R24 : label is "RVMAX";
ATTRIBUTE POWER of R24 : label is "RMAX";
ATTRIBUTE PSPICETEMPLATE of R24 : label is "R^@REFDES %1 %2 ?TOLERANCE|R^@REFDES| @VALUE TC=@TC1,@TC2 ?TOLERANCE|\n.model R^@REFDES RES R=1 DEV=@TOLERANCE% TC1=@TC1 TC2=@TC2|";


-- GATE INSTANCES

BEGIN
R25 : \1k\	PORT MAP(
	\2\ => N98425, 
	\1\ => N98451
);
R26 : \400\	PORT MAP(
	\2\ => N98201, 
	\1\ => GND
);
R27 : \50k\	PORT MAP(
	\2\ => N98633, 
	\1\ => N98621, 
	t => N98621
);
R28 : \50k\	PORT MAP(
	\2\ => N98691, 
	\1\ => GND, 
	t => GND
);
R29 : \10\	PORT MAP(
	\2\ => N98131, 
	\1\ => N98691
);
Q20 : QBC846B	PORT MAP(
	B => N98141, 
	E => N98233, 
	C => N97835
);
Q21 : QBC856B	PORT MAP(
	B => N97875, 
	E => N97965, 
	C => N97649
);
Q22 : QBC846B	PORT MAP(
	B => N97939, 
	E => N983391, 
	C => N97939
);
Q23 : QBC846B	PORT MAP(
	B => N97939, 
	E => N98425, 
	C => N98233
);
R30 : \10\	PORT MAP(
	\2\ => N98131, 
	\1\ => N98621
);
R31 : \200\	PORT MAP(
	\2\ => N97965, 
	\1\ => N97969
);
R32 : \50k\	PORT MAP(
	\2\ => N98201, 
	\1\ => N97983, 
	t => N97983
);
R33 : \1k\	PORT MAP(
	\2\ => N97649, 
	\1\ => N97755
);
TP2 : \V-\	PORT MAP(
	\1\ => N98451
);
R7 : \1k\	PORT MAP(
	\2\ => N98141, 
	\1\ => GND
);
TP3 : \TEST POINT\	PORT MAP(
	\1\ => N97755
);
R8 : \2k\	PORT MAP(
	\2\ => N98141, 
	\1\ => N97969
);
C6 : \33n\	PORT MAP(
	\1\ => N98633, 
	\2\ => N97965
);
C7 : \4.7u\	PORT MAP(
	\1\ => N97965, 
	\2\ => N97983
);
C8 : \33n\	PORT MAP(
	\1\ => GND, 
	\2\ => N98131
);
J1 : CON2	PORT MAP(
	\1\ => N97649, 
	\2\ => GND
);
J2 : CON2	PORT MAP(
	\1\ => N98451, 
	\2\ => GND
);
J3 : CON2	PORT MAP(
	\1\ => N98201, 
	\2\ => GND
);
D1 : D1N4148	PORT MAP(
	\1\ => N97969, 
	\2\ => N97965
);
R19 : \200\	PORT MAP(
	\2\ => N97649, 
	\1\ => N977031
);
D2 : D1N4148	PORT MAP(
	\1\ => N97965, 
	\2\ => N97969
);
D3 : \5V,LED,LED\	PORT MAP(
	\1\ => N97755, 
	\2\ => GND
);
Q17 : QBC856B	PORT MAP(
	B => N97835, 
	E => N977031, 
	C => N97875
);
Q18 : QBC856B	PORT MAP(
	B => N97835, 
	E => N977231, 
	C => N97835
);
Q19 : QBC846B	PORT MAP(
	B => N98131, 
	E => N98233, 
	C => N97875
);
R20 : \200\	PORT MAP(
	\2\ => N97649, 
	\1\ => N977231
);
R22 : \10k\	PORT MAP(
	\2\ => N97965, 
	\1\ => N98451
);
R23 : \4.7k\	PORT MAP(
	\2\ => N97649, 
	\1\ => N97939
);
R24 : \1k\	PORT MAP(
	\2\ => N983391, 
	\1\ => N98451
);
END STRUCTURE;

