-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Wednesday, December 03, 2025 14:49:36 GTB Standard Time

